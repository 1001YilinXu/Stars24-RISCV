//top.sv