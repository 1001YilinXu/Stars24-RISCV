package risc_pkg;
	parameter WORD_W = 32;
endpackage